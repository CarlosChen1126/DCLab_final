module DE2_115 (
	input CLOCK_50,
	input CLOCK2_50,
	input CLOCK3_50,
	input ENETCLK_25,
	input SMA_CLKIN,
	output SMA_CLKOUT,
	output [8:0] LEDG,
	output [17:0] LEDR,
	input [3:0] KEY,
	input [17:0] SW,
	output [6:0] HEX0,
	output [6:0] HEX1,
	output [6:0] HEX2,
	output [6:0] HEX3,
	output [6:0] HEX4,
	output [6:0] HEX5,
	output [6:0] HEX6,
	output [6:0] HEX7,
	output LCD_BLON,
	inout [7:0] LCD_DATA,
	output LCD_EN,
	output LCD_ON,
	output LCD_RS,
	output LCD_RW,
	output UART_CTS,
	input UART_RTS,
	input UART_RXD,
	output UART_TXD,
	inout PS2_CLK,
	inout PS2_DAT,
	inout PS2_CLK2,
	inout PS2_DAT2,
	output SD_CLK,
	inout SD_CMD,
	inout [3:0] SD_DAT,
	input SD_WP_N,
	output [7:0] VGA_B,
	output VGA_BLANK_N,
	output VGA_CLK,
	output [7:0] VGA_G,
	output VGA_HS,
	output [7:0] VGA_R,
	output VGA_SYNC_N,
	output VGA_VS,
	input AUD_ADCDAT,
	inout AUD_ADCLRCK,
	inout AUD_BCLK,
	output AUD_DACDAT,
	inout AUD_DACLRCK,
	output AUD_XCK,
	output EEP_I2C_SCLK,
	inout EEP_I2C_SDAT,
	output I2C_SCLK,
	inout I2C_SDAT,
	output ENET0_GTX_CLK,
	input ENET0_INT_N,
	output ENET0_MDC,
	input ENET0_MDIO,
	output ENET0_RST_N,
	input ENET0_RX_CLK,
	input ENET0_RX_COL,
	input ENET0_RX_CRS,
	input [3:0] ENET0_RX_DATA,
	input ENET0_RX_DV,
	input ENET0_RX_ER,
	input ENET0_TX_CLK,
	output [3:0] ENET0_TX_DATA,
	output ENET0_TX_EN,
	output ENET0_TX_ER,
	input ENET0_LINK100,
	output ENET1_GTX_CLK,
	input ENET1_INT_N,
	output ENET1_MDC,
	input ENET1_MDIO,
	output ENET1_RST_N,
	input ENET1_RX_CLK,
	input ENET1_RX_COL,
	input ENET1_RX_CRS,
	input [3:0] ENET1_RX_DATA,
	input ENET1_RX_DV,
	input ENET1_RX_ER,
	input ENET1_TX_CLK,
	output [3:0] ENET1_TX_DATA,
	output ENET1_TX_EN,
	output ENET1_TX_ER,
	input ENET1_LINK100,
	input TD_CLK27,
	input [7:0] TD_DATA,
	input TD_HS,
	output TD_RESET_N,
	input TD_VS,
	inout [15:0] OTG_DATA,
	output [1:0] OTG_ADDR,
	output OTG_CS_N,
	output OTG_WR_N,
	output OTG_RD_N,
	input OTG_INT,
	output OTG_RST_N,
	input IRDA_RXD,
	output [12:0] DRAM_ADDR,
	output [1:0] DRAM_BA,
	output DRAM_CAS_N,
	output DRAM_CKE,
	output DRAM_CLK,
	output DRAM_CS_N,
	inout [31:0] DRAM_DQ,
	output [3:0] DRAM_DQM,
	output DRAM_RAS_N,
	output DRAM_WE_N,
	output [19:0] SRAM_ADDR,
	output SRAM_CE_N,
	inout [15:0] SRAM_DQ,
	output SRAM_LB_N,
	output SRAM_OE_N,
	output SRAM_UB_N,
	output SRAM_WE_N,
	output [22:0] FL_ADDR,
	output FL_CE_N,
	inout [7:0] FL_DQ,
	output FL_OE_N,
	output FL_RST_N,
	input FL_RY,
	output FL_WE_N,
	output FL_WP_N,
	inout [35:0] GPIO,
	input HSMC_CLKIN_P1,
	input HSMC_CLKIN_P2,
	input HSMC_CLKIN0,
	output HSMC_CLKOUT_P1,
	output HSMC_CLKOUT_P2,
	output HSMC_CLKOUT0,
	inout [3:0] HSMC_D,
	input [16:0] HSMC_RX_D_P,
	output [16:0] HSMC_TX_D_P,
	inout [6:0] EX_IO
);

logic keydown_0,keydown_1,keydown_2;
logic CLK_25M, CLK_12M, CLK_100K;
logic [3:0] record;
logic [5:0] recd_time;


assign GPIO[9] = (state==3'd5);
assign AUD_XCK = CLK_12M;

vga_qsys qsys0(
	.clk_clk(CLOCK_50), 
	.reset_reset_n(KEY[3]),
	.clk100k_clk(CLK_100K),
	.clk25m_clk(CLK_25M),
	.clk12m_clk(CLK_12M)
);

Debounce deb0(
	.i_in(KEY[0]),
	.i_rst_n(KEY[3]),
	.i_clk(CLK_25M),
	.o_neg(keydown_0)
);
Debounce deb1(
	.i_in(KEY[1]),
	.i_rst_n(KEY[3]),
	.i_clk(CLK_25M),
	.o_neg(keydown_1)
);
logic music_in, music_stop;
Debounce deb2(
	.i_in(music_in),
	.i_rst_n(KEY[3]),
	.i_clk(CLK_12M),
	.o_neg(keydown_2)
);
logic [2:0] state;
logic [3:0] aud_state;
logic [1:0] music_index;
Top top0(
	.i_clk(CLOCK_50),
	.i_clk_25(CLK_25M),
	.i_rst_n(KEY[3]),
	.detect(GPIO[0]),
	.i_pos(GPIO[3:1]),
	.o_angle(GPIO[7:5]),
	.i_music_stop(music_stop),
	.VGA_R(VGA_R), 
	.VGA_G(VGA_G), 
	.VGA_B(VGA_B), 
	.VGA_CLK(VGA_CLK), 
	.VGA_BLANK_N(VGA_BLANK_N), 
	.VGA_HS(VGA_HS), 
	.VGA_VS(VGA_VS), 
	.VGA_SYNC_N(VGA_SYNC_N),
	.i_next(keydown_0),
	.i_finish_key(keydown_1),
	.state(state),
	.music_ind(music_index),
	.play_music(music_in)
);
logic [3:0] o_random_out;
Lfsr Lfsr0(
   .i_clk(CLK_12M),
   .i_rst_n(KEY[3]),
	.state(state),
   .o_random_out(o_random_out)
);
AudTop AudTop0(
	.i_rst_n(KEY[3]),
	.i_clk(CLK_12M),
	.i_key_0(keydown_2),
	.i_key_1(0),
	.i_key_2(0),
	.addr(addr),
	
	.music_stop(music_stop),
	
	.state(aud_state),
	
	// AudDSP and SRAM
	.i_speed({1'b0, o_random_out}), // design how user can decide mode on your own
	.i_fast(1),
	.i_slow_0(0),
	.i_slow_1(0),
	.sound_index(music_index),
	// AudDSP and SRAM
	.o_SRAM_ADDR(SRAM_ADDR), // [19:0]
	.io_SRAM_DQ(SRAM_DQ), 	 // [15:0]
	.o_SRAM_WE_N(SRAM_WE_N),
	.o_SRAM_CE_N(SRAM_CE_N),
	.o_SRAM_OE_N(SRAM_OE_N),
	.o_SRAM_LB_N(SRAM_LB_N),
	.o_SRAM_UB_N(SRAM_UB_N),
	
	// I2C
	.i_clk_100k(CLK_100K),
	.o_I2C_SCLK(I2C_SCLK),
	.io_I2C_SDAT(I2C_SDAT),
	
	// AudPlayer
	.i_AUD_ADCDAT(AUD_ADCDAT),
	.i_AUD_ADCLRCK(AUD_ADCLRCK),
	.i_AUD_BCLK(AUD_BCLK),
	.i_AUD_DACLRCK(AUD_DACLRCK),
	.o_AUD_DACDAT(AUD_DACDAT),

	// SEVENDECODER (optional display)
	.o_record_time(recd_time)
);
logic [19:0] addr;
SevenHexDecoder seven_dec0(
	.i_hex({1'b0,state}),
	.o_seven(HEX0)
);
SevenHexDecoder seven_dec1(
	.i_hex({3'd0,GPIO[0]}),
	.o_seven(HEX1)
);
SevenHexDecoder seven_dec2(
	.i_hex(addr[3:0]),
	.o_seven(HEX3)
);
SevenHexDecoder seven_dec3(
	.i_hex(addr[7:4]),
	.o_seven(HEX4)
);
SevenHexDecoder seven_dec4(
	.i_hex(addr[11:8]),
	.o_seven(HEX5)
);
//SevenHexDecoder seven_dec5(
//	.i_hex(addr[15:12]),
//	.o_seven(HEX6)
//);
//SevenHexDecoder seven_dec6(
//	.i_hex(addr[19:16]),
//	.o_seven(HEX7)
//);
SevenHexDecoder seven_dec5(
	.i_hex({1'b0,GPIO[7:5]}),
	.o_seven(HEX6)
);
SevenHexDecoder seven_dec6(
	.i_hex({1'b0,GPIO[3:1]}),
	.o_seven(HEX7)
);

//assign HEX1 = '1;
//assign HEX2 = '1;
//assign HEX3 = '1;
//assign HEX4 = '1;
//assign HEX5 = '1;
//assign HEX6 = '1;
//assign HEX7 = '1;

endmodule